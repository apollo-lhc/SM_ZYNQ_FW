default_top.vhd
--======================================================================
-- This may all look a bit cumbersome but in the context of ipbb and
-- friends it all works out quite well.
--======================================================================

use work.tcds2_interface_pkg.all;

package tcds2_interface_choice_mgt is

  constant C_TCDS2_BACKEND_MGT_TYPE : mgt_type_t := MGT_TYPE_GTHE4;

end package;

--======================================================================

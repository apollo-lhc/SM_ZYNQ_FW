module gf_add_5(op1, op2, res);

// -------------------------------------------------------------------------- //
// ------------- Triple Modular Redundancy Generator Directives ------------- //
// -------------------------------------------------------------------------- //
// tmrg do_not_touch
// -------------------------------------------------------------------------- //

	input      [4:0] op1; 
	input      [4:0] op2; 
	output     [4:0] res;

	assign res = op1 ^ op2;

endmodule

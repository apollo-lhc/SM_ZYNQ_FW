--====================================================================
-- Simply the choice of TCDS2 link medium: optical or electrical.
--====================================================================

package tcds2_link_medium_pkg is

  -- TCDS2 link medium: optical or electrical.
  type tcds2_link_medium_t is (TCDS2_LINK_MEDIUM_OPTICAL,
                               TCDS2_LINK_MEDIUM_ELECTRICAL);

end package;

--====================================================================

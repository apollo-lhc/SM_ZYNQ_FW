--======================================================================

use work.board_and_fw_id_pkg.all;

package constants_tcds2 is

  -- System ID: 'TCDS2'.
  constant c_SYSTEM_ID_TCDS2 : tcds2_id := "TCDS2   ";

  ----------

  -- The width of an IPBus word.
  constant C_IPBUS_WORD_WIDTH : integer := 32;

end constants_tcds2;

--======================================================================

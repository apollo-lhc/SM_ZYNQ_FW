library ieee;
use ieee.std_logic_1164.all;

use work.types.all;

entity SGMII_SI_data is
  
  port (
    entry : in  integer;
    addr  : out slv_12_t;
    data  : out slv_8_t);

end entity SGMII_SI_data;

architecture behavioral of SGMII_SI_data is

  --Upper 12  bits are addr, lower 12 are data
  constant writes : slv20_array_t(0 to 464) := (x"0B24C0",
                                                x"0B2500",
                                                x"054001",
                                                x"000600",
                                                x"000700",
                                                x"000800",
                                                x"000B68",
                                                x"001602",
                                                x"0017DC",
                                                x"0018EE",
                                                x"0019DD",
                                                x"001ADF",
                                                x"002B02",
                                                x"002C01",
                                                x"002D01",
                                                x"002E38",
                                                x"002F00",
                                                x"003000",
                                                x"003100",
                                                x"003200",
                                                x"003300",
                                                x"003400",
                                                x"003500",
                                                x"003638",
                                                x"003700",
                                                x"003800",
                                                x"003900",
                                                x"003A00",
                                                x"003B00",
                                                x"003C00",
                                                x"003D00",
                                                x"003F11",
                                                x"004004",
                                                x"00410D",
                                                x"004200",
                                                x"004300",
                                                x"004400",
                                                x"00450C",
                                                x"004632",
                                                x"004700",
                                                x"004800",
                                                x"004900",
                                                x"004A32",
                                                x"004B00",
                                                x"004C00",
                                                x"004D00",
                                                x"004E05",
                                                x"004F00",
                                                x"00500F",
                                                x"005103",
                                                x"005200",
                                                x"005300",
                                                x"005400",
                                                x"005503",
                                                x"005600",
                                                x"005700",
                                                x"005800",
                                                x"005901",
                                                x"005AAA",
                                                x"005BAA",
                                                x"005C0A",
                                                x"005D01",
                                                x"005E00",
                                                x"005F00",
                                                x"006000",
                                                x"006100",
                                                x"006200",
                                                x"006300",
                                                x"006400",
                                                x"006500",
                                                x"006600",
                                                x"006700",
                                                x"006800",
                                                x"006900",
                                                x"009202",
                                                x"0093A0",
                                                x"009500",
                                                x"009680",
                                                x"009860",
                                                x"009A02",
                                                x"009B60",
                                                x"009D08",
                                                x"009E40",
                                                x"00A020",
                                                x"00A200",
                                                x"00A9A7",
                                                x"00AA61",
                                                x"00AB00",
                                                x"00AC00",
                                                x"00E521",
                                                x"00EA0A",
                                                x"00EB60",
                                                x"00EC00",
                                                x"00ED00",
                                                x"010201",
                                                x"011202",
                                                x"011309",
                                                x"011433",
                                                x"011508",
                                                x"011702",
                                                x"011809",
                                                x"011933",
                                                x"011A08",
                                                x"012602",
                                                x"012709",
                                                x"012833",
                                                x"012909",
                                                x"012B02",
                                                x"012C09",
                                                x"012D33",
                                                x"012E0A",
                                                x"013F00",
                                                x"014000",
                                                x"014140",
                                                x"0142FF",
                                                x"020600",
                                                x"020832",
                                                x"020900",
                                                x"020A00",
                                                x"020B00",
                                                x"020C00",
                                                x"020D00",
                                                x"020E01",
                                                x"020F00",
                                                x"021000",
                                                x"021100",
                                                x"021200",
                                                x"021300",
                                                x"021400",
                                                x"021500",
                                                x"021600",
                                                x"021700",
                                                x"021800",
                                                x"021900",
                                                x"021A00",
                                                x"021B00",
                                                x"021C00",
                                                x"021D00",
                                                x"021E00",
                                                x"021F00",
                                                x"022000",
                                                x"022100",
                                                x"022200",
                                                x"022300",
                                                x"022400",
                                                x"022500",
                                                x"022600",
                                                x"022700",
                                                x"022800",
                                                x"022900",
                                                x"022A00",
                                                x"022B00",
                                                x"022C00",
                                                x"022D00",
                                                x"022E00",
                                                x"022F00",
                                                x"02310B",
                                                x"02320B",
                                                x"02330B",
                                                x"02340B",
                                                x"023500",
                                                x"023600",
                                                x"023700",
                                                x"0238C0",
                                                x"0239DA",
                                                x"023A00",
                                                x"023B00",
                                                x"023C00",
                                                x"023D00",
                                                x"023EC0",
                                                x"025003",
                                                x"025100",
                                                x"025200",
                                                x"025304",
                                                x"025400",
                                                x"025500",
                                                x"025C02",
                                                x"025D00",
                                                x"025E00",
                                                x"025F02",
                                                x"026000",
                                                x"026100",
                                                x"026B41",
                                                x"026C50",
                                                x"026D4F",
                                                x"026E4C",
                                                x"026F4C",
                                                x"02704F",
                                                x"027153",
                                                x"02724D",
                                                x"028A00",
                                                x"028B00",
                                                x"028C00",
                                                x"028D00",
                                                x"028E00",
                                                x"028F00",
                                                x"029000",
                                                x"029100",
                                                x"0294B0",
                                                x"029602",
                                                x"029702",
                                                x"029902",
                                                x"029DFA",
                                                x"029E01",
                                                x"029F00",
                                                x"02A9CC",
                                                x"02AA04",
                                                x"02AB00",
                                                x"02B7FF",
                                                x"030200",
                                                x"030300",
                                                x"030400",
                                                x"030500",
                                                x"030607",
                                                x"030700",
                                                x"030800",
                                                x"030900",
                                                x"030A00",
                                                x"030B80",
                                                x"030C00",
                                                x"030D00",
                                                x"030E00",
                                                x"030FEC",
                                                x"031060",
                                                x"031121",
                                                x"031200",
                                                x"031300",
                                                x"0314B8",
                                                x"0315C6",
                                                x"031692",
                                                x"031700",
                                                x"031800",
                                                x"0319C0",
                                                x"031A49",
                                                x"031B6E",
                                                x"031C0A",
                                                x"031D00",
                                                x"031E00",
                                                x"031F8B",
                                                x"032077",
                                                x"0321B7",
                                                x"032200",
                                                x"032300",
                                                x"032400",
                                                x"032500",
                                                x"032600",
                                                x"032700",
                                                x"032800",
                                                x"032900",
                                                x"032A00",
                                                x"032B00",
                                                x"032C00",
                                                x"032D00",
                                                x"033800",
                                                x"03391F",
                                                x"033B00",
                                                x"033C00",
                                                x"033D00",
                                                x"033E00",
                                                x"033F00",
                                                x"034000",
                                                x"034100",
                                                x"034200",
                                                x"034300",
                                                x"034400",
                                                x"034500",
                                                x"034600",
                                                x"034700",
                                                x"034800",
                                                x"034900",
                                                x"034A00",
                                                x"034B00",
                                                x"034C00",
                                                x"034D00",
                                                x"034E00",
                                                x"034F00",
                                                x"035000",
                                                x"035100",
                                                x"035200",
                                                x"035900",
                                                x"035A00",
                                                x"035B00",
                                                x"035C00",
                                                x"035D00",
                                                x"035E00",
                                                x"035F00",
                                                x"036000",
                                                x"048700",
                                                x"050813",
                                                x"050922",
                                                x"050A0C",
                                                x"050B0B",
                                                x"050C07",
                                                x"050D3F",
                                                x"050E16",
                                                x"050F2A",
                                                x"051009",
                                                x"051108",
                                                x"051207",
                                                x"05133F",
                                                x"051500",
                                                x"051600",
                                                x"051700",
                                                x"051800",
                                                x"0519BC",
                                                x"051A02",
                                                x"051B00",
                                                x"051C00",
                                                x"051D00",
                                                x"051E00",
                                                x"051F80",
                                                x"05212B",
                                                x"052A01",
                                                x"052B01",
                                                x"052C87",
                                                x"052D03",
                                                x"052E19",
                                                x"052F19",
                                                x"053100",
                                                x"053242",
                                                x"053303",
                                                x"053400",
                                                x"053500",
                                                x"053604",
                                                x"053700",
                                                x"053800",
                                                x"053900",
                                                x"053A02",
                                                x"053B03",
                                                x"053C00",
                                                x"053D11",
                                                x"053E06",
                                                x"05890D",
                                                x"058A00",
                                                x"059BFA",
                                                x"059D13",
                                                x"059E24",
                                                x"059F0C",
                                                x"05A00B",
                                                x"05A107",
                                                x"05A23F",
                                                x"05A603",
                                                x"080235",
                                                x"080305",
                                                x"080400",
                                                x"080500",
                                                x"080600",
                                                x"080700",
                                                x"080800",
                                                x"080900",
                                                x"080A00",
                                                x"080B00",
                                                x"080C00",
                                                x"080D00",
                                                x"080E00",
                                                x"080F00",
                                                x"081000",
                                                x"081100",
                                                x"081200",
                                                x"081300",
                                                x"081400",
                                                x"081500",
                                                x"081600",
                                                x"081700",
                                                x"081800",
                                                x"081900",
                                                x"081A00",
                                                x"081B00",
                                                x"081C00",
                                                x"081D00",
                                                x"081E00",
                                                x"081F00",
                                                x"082000",
                                                x"082100",
                                                x"082200",
                                                x"082300",
                                                x"082400",
                                                x"082500",
                                                x"082600",
                                                x"082700",
                                                x"082800",
                                                x"082900",
                                                x"082A00",
                                                x"082B00",
                                                x"082C00",
                                                x"082D00",
                                                x"082E00",
                                                x"082F00",
                                                x"083000",
                                                x"083100",
                                                x"083200",
                                                x"083300",
                                                x"083400",
                                                x"083500",
                                                x"083600",
                                                x"083700",
                                                x"083800",
                                                x"083900",
                                                x"083A00",
                                                x"083B00",
                                                x"083C00",
                                                x"083D00",
                                                x"083E00",
                                                x"083F00",
                                                x"084000",
                                                x"084100",
                                                x"084200",
                                                x"084300",
                                                x"084400",
                                                x"084500",
                                                x"084600",
                                                x"084700",
                                                x"084800",
                                                x"084900",
                                                x"084A00",
                                                x"084B00",
                                                x"084C00",
                                                x"084D00",
                                                x"084E00",
                                                x"084F00",
                                                x"085000",
                                                x"085100",
                                                x"085200",
                                                x"085300",
                                                x"085400",
                                                x"085500",
                                                x"085600",
                                                x"085700",
                                                x"085800",
                                                x"085900",
                                                x"085A00",
                                                x"085B00",
                                                x"085C00",
                                                x"085D00",
                                                x"085E00",
                                                x"085F00",
                                                x"086000",
                                                x"086100",
                                                x"090E02",
                                                x"094300",
                                                x"094901",
                                                x"094A01",
                                                x"094E49",
                                                x"094F02",
                                                x"095E00",
                                                x"0A0200",
                                                x"0A0307",
                                                x"0A0401",
                                                x"0A0507",
                                                x"0A1400",
                                                x"0A1A00",
                                                x"0A2000",
                                                x"0A2600",
                                                x"0B442F",
                                                x"0B4600",
                                                x"0B470E",
                                                x"0B480E",
                                                x"0B4A08",
                                                x"0B570E",
                                                x"0B5801",
                                                x"051401",
                                                x"001C01",
                                                x"054000",
                                                x"0B24C3",
                                                x"0B2502"
                                                );
--  constant writes : slv20_array_t(0 to 464) := (x"B24C0",
--                                              x"B2500",
--                                              x"54001",
--                                              x"00600",
--                                              x"00700",
--                                              x"00800",
--                                              x"00B68",
--                                              x"01602",
--                                              x"017DC",
--                                              x"018EE",
--                                              x"019DD",
--                                              x"01ADF",
--                                              x"02B02",
--                                              x"02C01",
--                                              x"02D01",
--                                              x"02E38",
--                                              x"02F00",
--                                              x"03000",
--                                              x"03100",
--                                              x"03200",
--                                              x"03300",
--                                              x"03400",
--                                              x"03500",
--                                              x"03638",
--                                              x"03700",
--                                              x"03800",
--                                              x"03900",
--                                              x"03A00",
--                                              x"03B00",
--                                              x"03C00",
--                                              x"03D00",
--                                              x"03F11",
--                                              x"04004",
--                                              x"0410D",
--                                              x"04200",
--                                              x"04300",
--                                              x"04400",
--                                              x"0450C",
--                                              x"04632",
--                                              x"04700",
--                                              x"04800",
--                                              x"04900",
--                                              x"04A32",
--                                              x"04B00",
--                                              x"04C00",
--                                              x"04D00",
--                                              x"04E05",
--                                              x"04F00",
--                                              x"0500F",
--                                              x"05103",
--                                              x"05200",
--                                              x"05300",
--                                              x"05400",
--                                              x"05503",
--                                              x"05600",
--                                              x"05700",
--                                              x"05800",
--                                              x"05901",
--                                              x"05AAA",
--                                              x"05BAA",
--                                              x"05C0A",
--                                              x"05D01",
--                                              x"05E00",
--                                              x"05F00",
--                                              x"06000",
--                                              x"06100",
--                                              x"06200",
--                                              x"06300",
--                                              x"06400",
--                                              x"06500",
--                                              x"06600",
--                                              x"06700",
--                                              x"06800",
--                                              x"06900",
--                                              x"09202",
--                                              x"093A0",
--                                              x"09500",
--                                              x"09680",
--                                              x"09860",
--                                              x"09A02",
--                                              x"09B60",
--                                              x"09D08",
--                                              x"09E40",
--                                              x"0A020",
--                                              x"0A200",
--                                              x"0A9A7",
--                                              x"0AA61",
--                                              x"0AB00",
--                                              x"0AC00",
--                                              x"0E521",
--                                              x"0EA0A",
--                                              x"0EB60",
--                                              x"0EC00",
--                                              x"0ED00",
--                                              x"10201",
--                                              x"11202",
--                                              x"11309",
--                                              x"11433",
--                                              x"11508",
--                                              x"11702",
--                                              x"11809",
--                                              x"11933",
--                                              x"11A08",
--                                              x"12602",
--                                              x"12709",
--                                              x"12833",
--                                              x"12909",
--                                              x"12B02",
--                                              x"12C09",
--                                              x"12D33",
--                                              x"12E0A",
--                                              x"13F00",
--                                              x"14000",
--                                              x"14140",
--                                              x"142FF",
--                                              x"20600",
--                                              x"20832",
--                                              x"20900",
--                                              x"20A00",
--                                              x"20B00",
--                                              x"20C00",
--                                              x"20D00",
--                                              x"20E01",
--                                              x"20F00",
--                                              x"21000",
--                                              x"21100",
--                                              x"21200",
--                                              x"21300",
--                                              x"21400",
--                                              x"21500",
--                                              x"21600",
--                                              x"21700",
--                                              x"21800",
--                                              x"21900",
--                                              x"21A00",
--                                              x"21B00",
--                                              x"21C00",
--                                              x"21D00",
--                                              x"21E00",
--                                              x"21F00",
--                                              x"22000",
--                                              x"22100",
--                                              x"22200",
--                                              x"22300",
--                                              x"22400",
--                                              x"22500",
--                                              x"22600",
--                                              x"22700",
--                                              x"22800",
--                                              x"22900",
--                                              x"22A00",
--                                              x"22B00",
--                                              x"22C00",
--                                              x"22D00",
--                                              x"22E00",
--                                              x"22F00",
--                                              x"2310B",
--                                              x"2320B",
--                                              x"2330B",
--                                              x"2340B",
--                                              x"23500",
--                                              x"23600",
--                                              x"23700",
--                                              x"238C0",
--                                              x"239DA",
--                                              x"23A00",
--                                              x"23B00",
--                                              x"23C00",
--                                              x"23D00",
--                                              x"23EC0",
--                                              x"25003",
--                                              x"25100",
--                                              x"25200",
--                                              x"25304",
--                                              x"25400",
--                                              x"25500",
--                                              x"25C02",
--                                              x"25D00",
--                                              x"25E00",
--                                              x"25F02",
--                                              x"26000",
--                                              x"26100",
--                                              x"26B41",
--                                              x"26C50",
--                                              x"26D4F",
--                                              x"26E4C",
--                                              x"26F4C",
--                                              x"2704F",
--                                              x"27153",
--                                              x"2724D",
--                                              x"28A00",
--                                              x"28B00",
--                                              x"28C00",
--                                              x"28D00",
--                                              x"28E00",
--                                              x"28F00",
--                                              x"29000",
--                                              x"29100",
--                                              x"294B0",
--                                              x"29602",
--                                              x"29702",
--                                              x"29902",
--                                              x"29DFA",
--                                              x"29E01",
--                                              x"29F00",
--                                              x"2A9CC",
--                                              x"2AA04",
--                                              x"2AB00",
--                                              x"2B7FF",
--                                              x"30200",
--                                              x"30300",
--                                              x"30400",
--                                              x"30500",
--                                              x"30607",
--                                              x"30700",
--                                              x"30800",
--                                              x"30900",
--                                              x"30A00",
--                                              x"30B80",
--                                              x"30C00",
--                                              x"30D00",
--                                              x"30E00",
--                                              x"30FEC",
--                                              x"31060",
--                                              x"31121",
--                                              x"31200",
--                                              x"31300",
--                                              x"314B8",
--                                              x"315C6",
--                                              x"31692",
--                                              x"31700",
--                                              x"31800",
--                                              x"319C0",
--                                              x"31A49",
--                                              x"31B6E",
--                                              x"31C0A",
--                                              x"31D00",
--                                              x"31E00",
--                                              x"31F8B",
--                                              x"32077",
--                                              x"321B7",
--                                              x"32200",
--                                              x"32300",
--                                              x"32400",
--                                              x"32500",
--                                              x"32600",
--                                              x"32700",
--                                              x"32800",
--                                              x"32900",
--                                              x"32A00",
--                                              x"32B00",
--                                              x"32C00",
--                                              x"32D00",
--                                              x"33800",
--                                              x"3391F",
--                                              x"33B00",
--                                              x"33C00",
--                                              x"33D00",
--                                              x"33E00",
--                                              x"33F00",
--                                              x"34000",
--                                              x"34100",
--                                              x"34200",
--                                              x"34300",
--                                              x"34400",
--                                              x"34500",
--                                              x"34600",
--                                              x"34700",
--                                              x"34800",
--                                              x"34900",
--                                              x"34A00",
--                                              x"34B00",
--                                              x"34C00",
--                                              x"34D00",
--                                              x"34E00",
--                                              x"34F00",
--                                              x"35000",
--                                              x"35100",
--                                              x"35200",
--                                              x"35900",
--                                              x"35A00",
--                                              x"35B00",
--                                              x"35C00",
--                                              x"35D00",
--                                              x"35E00",
--                                              x"35F00",
--                                              x"36000",
--                                              x"48700",
--                                              x"50813",
--                                              x"50922",
--                                              x"50A0C",
--                                              x"50B0B",
--                                              x"50C07",
--                                              x"50D3F",
--                                              x"50E16",
--                                              x"50F2A",
--                                              x"51009",
--                                              x"51108",
--                                              x"51207",
--                                              x"5133F",
--                                              x"51500",
--                                              x"51600",
--                                              x"51700",
--                                              x"51800",
--                                              x"519BC",
--                                              x"51A02",
--                                              x"51B00",
--                                              x"51C00",
--                                              x"51D00",
--                                              x"51E00",
--                                              x"51F80",
--                                              x"5212B",
--                                              x"52A01",
--                                              x"52B01",
--                                              x"52C87",
--                                              x"52D03",
--                                              x"52E19",
--                                              x"52F19",
--                                              x"53100",
--                                              x"53242",
--                                              x"53303",
--                                              x"53400",
--                                              x"53500",
--                                              x"53604",
--                                              x"53700",
--                                              x"53800",
--                                              x"53900",
--                                              x"53A02",
--                                              x"53B03",
--                                              x"53C00",
--                                              x"53D11",
--                                              x"53E06",
--                                              x"5890D",
--                                              x"58A00",
--                                              x"59BFA",
--                                              x"59D13",
--                                              x"59E24",
--                                              x"59F0C",
--                                              x"5A00B",
--                                              x"5A107",
--                                              x"5A23F",
--                                              x"5A603",
--                                              x"80235",
--                                              x"80305",
--                                              x"80400",
--                                              x"80500",
--                                              x"80600",
--                                              x"80700",
--                                              x"80800",
--                                              x"80900",
--                                              x"80A00",
--                                              x"80B00",
--                                              x"80C00",
--                                              x"80D00",
--                                              x"80E00",
--                                              x"80F00",
--                                              x"81000",
--                                              x"81100",
--                                              x"81200",
--                                              x"81300",
--                                              x"81400",
--                                              x"81500",
--                                              x"81600",
--                                              x"81700",
--                                              x"81800",
--                                              x"81900",
--                                              x"81A00",
--                                              x"81B00",
--                                              x"81C00",
--                                              x"81D00",
--                                              x"81E00",
--                                              x"81F00",
--                                              x"82000",
--                                              x"82100",
--                                              x"82200",
--                                              x"82300",
--                                              x"82400",
--                                              x"82500",
--                                              x"82600",
--                                              x"82700",
--                                              x"82800",
--                                              x"82900",
--                                              x"82A00",
--                                              x"82B00",
--                                              x"82C00",
--                                              x"82D00",
--                                              x"82E00",
--                                              x"82F00",
--                                              x"83000",
--                                              x"83100",
--                                              x"83200",
--                                              x"83300",
--                                              x"83400",
--                                              x"83500",
--                                              x"83600",
--                                              x"83700",
--                                              x"83800",
--                                              x"83900",
--                                              x"83A00",
--                                              x"83B00",
--                                              x"83C00",
--                                              x"83D00",
--                                              x"83E00",
--                                              x"83F00",
--                                              x"84000",
--                                              x"84100",
--                                              x"84200",
--                                              x"84300",
--                                              x"84400",
--                                              x"84500",
--                                              x"84600",
--                                              x"84700",
--                                              x"84800",
--                                              x"84900",
--                                              x"84A00",
--                                              x"84B00",
--                                              x"84C00",
--                                              x"84D00",
--                                              x"84E00",
--                                              x"84F00",
--                                              x"85000",
--                                              x"85100",
--                                              x"85200",
--                                              x"85300",
--                                              x"85400",
--                                              x"85500",
--                                              x"85600",
--                                              x"85700",
--                                              x"85800",
--                                              x"85900",
--                                              x"85A00",
--                                              x"85B00",
--                                              x"85C00",
--                                              x"85D00",
--                                              x"85E00",
--                                              x"85F00",
--                                              x"86000",
--                                              x"86100",
--                                              x"90E02",
--                                              x"94300",
--                                              x"94901",
--                                              x"94A01",
--                                              x"94E49",
--                                              x"94F02",
--                                              x"95E00",
--                                              x"A0200",
--                                              x"A0307",
--                                              x"A0401",
--                                              x"A0507",
--                                              x"A1400",
--                                              x"A1A00",
--                                              x"A2000",
--                                              x"A2600",
--                                              x"B442F",
--                                              x"B4600",
--                                              x"B470E",
--                                              x"B480E",
--                                              x"B4A08",
--                                              x"B570E",
--                                              x"B5801",
--                                              x"51401",
--                                              x"01C01",
--                                              x"54000",
--                                              x"B24C3",
--                                              x"B2502"
--                                              );
begin  -- architecture behavioral

  addr <= writes(entry)(19 downto 8);
  data <= writes(entry)( 7 downto 0);

end architecture behavioral;

../rev2_xc7z035/src/top.vhd
top_rev2_xc7z035.vhd
------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : lhc_support.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module LHC_support
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
--***********************************Entity Declaration************************

entity LHC_support is
  generic
    (
      EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
      STABLE_CLOCK_PERIOD                     : integer   := 16  

      );
  port
    (
      SOFT_RESET_TX_IN                        : in   std_logic;
      SOFT_RESET_RX_IN                        : in   std_logic;
      DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;

      GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
      GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
      GT0_DATA_VALID_IN                       : in   std_logic;
      GT0_TX_MMCM_LOCK_OUT                    : out  std_logic;
      GT0_RX_MMCM_LOCK_OUT                    : out  std_logic;
      
      GT0_TXUSRCLK_OUT                        : out  std_logic;
      GT0_TXUSRCLK2_OUT                       : out  std_logic;
      GT0_RXUSRCLK_OUT                        : out  std_logic;
      GT0_RXUSRCLK2_OUT                       : out  std_logic;

      --_________________________________________________________________________
      --GT0  (X1Y13)
      --____________________________CHANNEL PORTS________________________________
      --------------------------------- CPLL Ports -------------------------------
      gt0_cpllfbclklost_out                   : out  std_logic;
      gt0_cplllock_out                        : out  std_logic;
      gt0_cpllreset_in                        : in   std_logic;
      ---------------------------- Channel - DRP Ports  --------------------------
      gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
      gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
      gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
      gt0_drpen_in                            : in   std_logic;
      gt0_drprdy_out                          : out  std_logic;
      gt0_drpwe_in                            : in   std_logic;
      --------------------------- Digital Monitor Ports --------------------------
      gt0_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
      --------------------- RX Initialization and Reset Ports --------------------
      gt0_eyescanreset_in                     : in   std_logic;
      gt0_rxuserrdy_in                        : in   std_logic;
      -------------------------- RX Margin Analysis Ports ------------------------
      gt0_eyescandataerror_out                : out  std_logic;
      gt0_eyescantrigger_in                   : in   std_logic;
      ------------------ Receive Ports - FPGA RX interface Ports -----------------
      gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
      ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
      gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
      gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
      --------------------------- Receive Ports - RX AFE -------------------------
      gt0_gtxrxp_in                           : in   std_logic;
      ------------------------ Receive Ports - RX AFE Ports ----------------------
      gt0_gtxrxn_in                           : in   std_logic;
      --------------------- Receive Ports - RX Equalizer Ports -------------------
      gt0_rxdfelpmreset_in                    : in   std_logic;
      gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
      gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
      --------------- Receive Ports - RX Fabric Output Control Ports -------------
      gt0_rxoutclkfabric_out                  : out  std_logic;
      ------------- Receive Ports - RX Initialization and Reset Ports ------------
      gt0_gtrxreset_in                        : in   std_logic;
      gt0_rxpmareset_in                       : in   std_logic;
      ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
      gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
      -------------- Receive Ports -RX Initialization and Reset Ports ------------
      gt0_rxresetdone_out                     : out  std_logic;
      --------------------- TX Initialization and Reset Ports --------------------
      gt0_gttxreset_in                        : in   std_logic;
      gt0_txuserrdy_in                        : in   std_logic;
      ------------------ Transmit Ports - TX Data Path interface -----------------
      gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
      ---------------- Transmit Ports - TX Driver and OOB signaling --------------
      gt0_gtxtxn_out                          : out  std_logic;
      gt0_gtxtxp_out                          : out  std_logic;
      ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
      gt0_txoutclkfabric_out                  : out  std_logic;
      gt0_txoutclkpcs_out                     : out  std_logic;
      --------------------- Transmit Ports - TX Gearbox Ports --------------------
      gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
      ------------- Transmit Ports - TX Initialization and Reset Ports -----------
      gt0_txresetdone_out                     : out  std_logic;

      --____________________________COMMON PORTS________________________________
      GT0_QPLLOUTCLK_OUT    : in  std_logic;
      GT0_QPLLOUTREFCLK_OUT : in  std_logic;
      Q3_CLK1_GTREFCLK_OUT  : in  std_logic;
      sysclk_in             : in  std_logic

      );

end LHC_support;

architecture RTL of LHC_support is
  attribute DowngradeIPIdentifiedWarnings: string;
  attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

--**************************Component Declarations*****************************

  component LHC
    
    port
      (
        SYSCLK_IN                               : in   std_logic;
        SOFT_RESET_TX_IN                        : in   std_logic;
        SOFT_RESET_RX_IN                        : in   std_logic;
        DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
        GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
        GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
        GT0_DATA_VALID_IN                       : in   std_logic;
        GT0_TX_MMCM_LOCK_IN                     : in   std_logic;
        GT0_TX_MMCM_RESET_OUT                   : out  std_logic;
        GT0_RX_MMCM_LOCK_IN                     : in   std_logic;
        GT0_RX_MMCM_RESET_OUT                   : out  std_logic;

        --_________________________________________________________________________
        --GT0  (X1Y13)
        --____________________________CHANNEL PORTS________________________________
        --------------------------------- CPLL Ports -------------------------------
        gt0_cpllfbclklost_out                   : out  std_logic;
        gt0_cplllock_out                        : out  std_logic;
        gt0_cplllockdetclk_in                   : in   std_logic;
        gt0_cpllreset_in                        : in   std_logic;
        -------------------------- Channel - Clocking Ports ------------------------
        gt0_gtrefclk0_in                        : in   std_logic;
        gt0_gtrefclk1_in                        : in   std_logic;
        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
        gt0_drpclk_in                           : in   std_logic;
        gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
        gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
        gt0_drpen_in                            : in   std_logic;
        gt0_drprdy_out                          : out  std_logic;
        gt0_drpwe_in                            : in   std_logic;
        --------------------------- Digital Monitor Ports --------------------------
        gt0_dmonitorout_out                     : out  std_logic_vector(7 downto 0);
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in                     : in   std_logic;
        gt0_rxuserrdy_in                        : in   std_logic;
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out                : out  std_logic;
        gt0_eyescantrigger_in                   : in   std_logic;
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxusrclk_in                         : in   std_logic;
        gt0_rxusrclk2_in                        : in   std_logic;
        ------------------ Receive Ports - FPGA RX interface Ports -----------------
        gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
        gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
        --------------------------- Receive Ports - RX AFE -------------------------
        gt0_gtxrxp_in                           : in   std_logic;
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gtxrxn_in                           : in   std_logic;
        --------------------- Receive Ports - RX Equalizer Ports -------------------
        gt0_rxdfelpmreset_in                    : in   std_logic;
        gt0_rxmonitorout_out                    : out  std_logic_vector(6 downto 0);
        gt0_rxmonitorsel_in                     : in   std_logic_vector(1 downto 0);
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclkfabric_out                  : out  std_logic;
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                        : in   std_logic;
        gt0_rxpmareset_in                       : in   std_logic;
        ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
        gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out                     : out  std_logic;
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                        : in   std_logic;
        gt0_txuserrdy_in                        : in   std_logic;
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txusrclk_in                         : in   std_logic;
        gt0_txusrclk2_in                        : in   std_logic;
        ------------------ Transmit Ports - TX Data Path interface -----------------
        gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
        ---------------- Transmit Ports - TX Driver and OOB signaling --------------
        gt0_gtxtxn_out                          : out  std_logic;
        gt0_gtxtxp_out                          : out  std_logic;
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                        : out  std_logic;
        gt0_txoutclkfabric_out                  : out  std_logic;
        gt0_txoutclkpcs_out                     : out  std_logic;
        --------------------- Transmit Ports - TX Gearbox Ports --------------------
        gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out                     : out  std_logic;


        --____________________________COMMON PORTS________________________________
        GT0_QPLLOUTCLK_IN  : in std_logic;
        GT0_QPLLOUTREFCLK_IN : in std_logic

        );

  end component;

  component LHC_GT_USRCLK_SOURCE 
    port
      (
        
        GT0_TXUSRCLK_OUT             : out std_logic;
        GT0_TXUSRCLK2_OUT            : out std_logic;
        GT0_TXOUTCLK_IN              : in  std_logic;
        GT0_TXCLK_LOCK_OUT           : out std_logic;
        GT0_TX_MMCM_RESET_IN         : in std_logic;
        GT0_RXUSRCLK_OUT             : out std_logic;
        GT0_RXUSRCLK2_OUT            : out std_logic;
        GT0_RXCLK_LOCK_OUT           : out std_logic;
        GT0_RX_MMCM_RESET_IN         : in std_logic
        );
  end component;

--***********************************Parameter Declarations********************

  constant DLY : time := 1 ns;

--************************** Register Declarations ****************************

  signal   gt0_txfsmresetdone_i            : std_logic;
  signal   gt0_rxfsmresetdone_i            : std_logic;
  signal   gt0_txfsmresetdone_r            : std_logic;
  signal   gt0_txfsmresetdone_r2           : std_logic;
  signal   gt0_rxresetdone_r               : std_logic;
  signal   gt0_rxresetdone_r2              : std_logic;
  signal   gt0_rxresetdone_r3              : std_logic;


  signal   reset_pulse                     : std_logic_vector(3 downto 0);
  signal   reset_counter  :   unsigned(5 downto 0) := "000000";

--**************************** Wire Declarations ******************************
  -------------------------- GT Wrapper Wires ------------------------------
  --________________________________________________________________________
  --________________________________________________________________________
  --GT0  (X1Y13)

  --------------------------------- CPLL Ports -------------------------------
  signal  gt0_cpllfbclklost_i             : std_logic;
  signal  gt0_cplllock_i                  : std_logic;
  signal  gt0_cpllrefclklost_i            : std_logic;
  signal  gt0_cpllreset_i                 : std_logic;
  ---------------------------- Channel - DRP Ports  --------------------------
  signal  gt0_drpaddr_i                   : std_logic_vector(8 downto 0);
  signal  gt0_drpdi_i                     : std_logic_vector(15 downto 0);
  signal  gt0_drpdo_i                     : std_logic_vector(15 downto 0);
  signal  gt0_drpen_i                     : std_logic;
  signal  gt0_drprdy_i                    : std_logic;
  signal  gt0_drpwe_i                     : std_logic;
  --------------------------- Digital Monitor Ports --------------------------
  signal  gt0_dmonitorout_i               : std_logic_vector(7 downto 0);
  --------------------- RX Initialization and Reset Ports --------------------
  signal  gt0_eyescanreset_i              : std_logic;
  signal  gt0_rxuserrdy_i                 : std_logic;
  -------------------------- RX Margin Analysis Ports ------------------------
  signal  gt0_eyescandataerror_i          : std_logic;
  signal  gt0_eyescantrigger_i            : std_logic;
  ------------------ Receive Ports - FPGA RX interface Ports -----------------
  signal  gt0_rxdata_i                    : std_logic_vector(31 downto 0);
  ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
  signal  gt0_rxdisperr_i                 : std_logic_vector(3 downto 0);
  signal  gt0_rxnotintable_i              : std_logic_vector(3 downto 0);
  --------------------------- Receive Ports - RX AFE -------------------------
  signal  gt0_gtxrxp_i                    : std_logic;
  ------------------------ Receive Ports - RX AFE Ports ----------------------
  signal  gt0_gtxrxn_i                    : std_logic;
  -------------------- Receive Ports - RX Equailizer Ports -------------------
  signal  gt0_rxlpmhfhold_i               : std_logic;
  signal  gt0_rxlpmlfhold_i               : std_logic;
  --------------------- Receive Ports - RX Equalizer Ports -------------------
  signal  gt0_rxdfelpmreset_i             : std_logic;
  signal  gt0_rxmonitorout_i              : std_logic_vector(6 downto 0);
  signal  gt0_rxmonitorsel_i              : std_logic_vector(1 downto 0);
  --------------- Receive Ports - RX Fabric Output Control Ports -------------
  signal  gt0_rxoutclk_i                  : std_logic;
  signal  gt0_rxoutclkfabric_i            : std_logic;
  ------------- Receive Ports - RX Initialization and Reset Ports ------------
  signal  gt0_gtrxreset_i                 : std_logic;
  signal  gt0_rxpmareset_i                : std_logic;
  ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
  signal  gt0_rxcharisk_i                 : std_logic_vector(3 downto 0);
  -------------- Receive Ports -RX Initialization and Reset Ports ------------
  signal  gt0_rxresetdone_i               : std_logic;
  --------------------- TX Initialization and Reset Ports --------------------
  signal  gt0_gttxreset_i                 : std_logic;
  signal  gt0_txuserrdy_i                 : std_logic;
  ------------------ Transmit Ports - TX Data Path interface -----------------
  signal  gt0_txdata_i                    : std_logic_vector(31 downto 0);
  ---------------- Transmit Ports - TX Driver and OOB signaling --------------
  signal  gt0_gtxtxn_i                    : std_logic;
  signal  gt0_gtxtxp_i                    : std_logic;
  ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
  signal  gt0_txoutclk_i                  : std_logic;
  signal  gt0_txoutclkfabric_i            : std_logic;
  signal  gt0_txoutclkpcs_i               : std_logic;
  --------------------- Transmit Ports - TX Gearbox Ports --------------------
  signal  gt0_txcharisk_i                 : std_logic_vector(3 downto 0);
  ------------- Transmit Ports - TX Initialization and Reset Ports -----------
  signal  gt0_txresetdone_i               : std_logic;

  --____________________________COMMON PORTS________________________________
  signal gt0_qpllreset_i  : std_logic;

  ------------------------------- Global Signals -----------------------------
  signal  gt0_tx_system_reset_c           : std_logic;
  signal  gt0_rx_system_reset_c           : std_logic;
  signal  tied_to_ground_i                : std_logic;
  signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
  signal  tied_to_vcc_i                   : std_logic;
  signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
  signal  drpclk_in_i                     : std_logic;
  signal  sysclk_in_i                     : std_logic;
  signal  GTTXRESET_IN                    : std_logic;
  signal  GTRXRESET_IN                    : std_logic;
  signal  CPLLRESET_IN                    : std_logic;
  signal  QPLLRESET_IN                    : std_logic;

  attribute keep: string;
  ------------------------------- User Clocks ---------------------------------
  signal    gt0_txusrclk_i                  : std_logic; 
  signal    gt0_txusrclk2_i                 : std_logic; 
  signal    gt0_rxusrclk_i                  : std_logic; 
  signal    gt0_rxusrclk2_i                 : std_logic; 
  
  
  
  
  signal    gt0_txmmcm_lock_i               : std_logic;
  signal    gt0_txmmcm_reset_i              : std_logic;
  signal    gt0_rxmmcm_lock_i               : std_logic; 
  signal    gt0_rxmmcm_reset_i              : std_logic;
--**************************** Main Body of Code *******************************
begin

  --  Static signal Assigments
  tied_to_ground_i                             <= '0';
  tied_to_ground_vec_i                         <= x"0000000000000000";
  tied_to_vcc_i                                <= '1';
  tied_to_vcc_vec_i                            <= "11111111";

  GT0_TX_MMCM_LOCK_OUT <= gt0_txmmcm_lock_i;
  GT0_RX_MMCM_LOCK_OUT <= gt0_rxmmcm_lock_i;
  

  
  GT0_TXUSRCLK_OUT <= gt0_txusrclk_i; 
  GT0_TXUSRCLK2_OUT <= gt0_txusrclk2_i;
  GT0_RXUSRCLK_OUT <= gt0_rxusrclk_i;
  GT0_RXUSRCLK2_OUT <= gt0_rxusrclk2_i;


  
  
  gt_usrclk_source : LHC_GT_USRCLK_SOURCE
    port map
    (
      
      GT0_TXUSRCLK_OUT                =>      gt0_txusrclk_i,
      GT0_TXUSRCLK2_OUT               =>      gt0_txusrclk2_i,
      GT0_TXOUTCLK_IN                 =>      gt0_txoutclk_i,
      GT0_TXCLK_LOCK_OUT              =>      gt0_txmmcm_lock_i,
      GT0_TX_MMCM_RESET_IN            =>      gt0_txmmcm_reset_i,
      GT0_RXUSRCLK_OUT                =>      gt0_rxusrclk_i,
      GT0_RXUSRCLK2_OUT               =>      gt0_rxusrclk2_i,
      GT0_RXCLK_LOCK_OUT              =>      gt0_rxmmcm_lock_i,
      GT0_RX_MMCM_RESET_IN            =>      gt0_rxmmcm_reset_i
      );

  sysclk_in_i <= sysclk_in;


  LHC_init_i : LHC
    port map
    (
      sysclk_in                       =>      sysclk_in_i,
      soft_reset_tx_in                =>      SOFT_RESET_TX_IN,
      soft_reset_rx_in                =>      SOFT_RESET_RX_IN,
      dont_reset_on_data_error_in     =>      DONT_RESET_ON_DATA_ERROR_IN,
      gt0_tx_mmcm_lock_in             =>      gt0_txmmcm_lock_i,
      gt0_tx_mmcm_reset_out           =>      gt0_txmmcm_reset_i,
      gt0_rx_mmcm_lock_in             =>      gt0_rxmmcm_lock_i,
      gt0_rx_mmcm_reset_out           =>      gt0_rxmmcm_reset_i,
      gt0_tx_fsm_reset_done_out       =>      gt0_tx_fsm_reset_done_out,
      gt0_rx_fsm_reset_done_out       =>      gt0_rx_fsm_reset_done_out,
      gt0_data_valid_in               =>      gt0_data_valid_in,

      --_____________________________________________________________________
      --_____________________________________________________________________
      --GT0  (X1Y13)

      --------------------------------- CPLL Ports -------------------------------
      gt0_cpllfbclklost_out           =>      gt0_cpllfbclklost_out,
      gt0_cplllock_out                =>      gt0_cplllock_out,
      gt0_cplllockdetclk_in           =>      sysclk_in_i,
      gt0_cpllreset_in                =>      gt0_cpllreset_in,
      -------------------------- Channel - Clocking Ports ------------------------
      gt0_gtrefclk0_in                =>      tied_to_ground_i,
      gt0_gtrefclk1_in                =>      Q3_CLK1_GTREFCLK_OUT,
      ---------------------------- Channel - DRP Ports  --------------------------
      gt0_drpaddr_in                  =>      gt0_drpaddr_in,
      gt0_drpclk_in                   =>      sysclk_in_i,
      gt0_drpdi_in                    =>      gt0_drpdi_in,
      gt0_drpdo_out                   =>      gt0_drpdo_out,
      gt0_drpen_in                    =>      gt0_drpen_in,
      gt0_drprdy_out                  =>      gt0_drprdy_out,
      gt0_drpwe_in                    =>      gt0_drpwe_in,
      --------------------------- Digital Monitor Ports --------------------------
      gt0_dmonitorout_out             =>      gt0_dmonitorout_out,
      --------------------- RX Initialization and Reset Ports --------------------
      gt0_eyescanreset_in             =>      gt0_eyescanreset_in,
      gt0_rxuserrdy_in                =>      gt0_rxuserrdy_in,
      -------------------------- RX Margin Analysis Ports ------------------------
      gt0_eyescandataerror_out        =>      gt0_eyescandataerror_out,
      gt0_eyescantrigger_in           =>      gt0_eyescantrigger_in,
      ------------------ Receive Ports - FPGA RX Interface Ports -----------------
      gt0_rxusrclk_in                 =>      gt0_rxusrclk_i,
      gt0_rxusrclk2_in                =>      gt0_rxusrclk2_i,
      ------------------ Receive Ports - FPGA RX interface Ports -----------------
      gt0_rxdata_out                  =>      gt0_rxdata_out,
      ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
      gt0_rxdisperr_out               =>      gt0_rxdisperr_out,
      gt0_rxnotintable_out            =>      gt0_rxnotintable_out,
      --------------------------- Receive Ports - RX AFE -------------------------
      gt0_gtxrxp_in                   =>      gt0_gtxrxp_in,
      ------------------------ Receive Ports - RX AFE Ports ----------------------
      gt0_gtxrxn_in                   =>      gt0_gtxrxn_in,
      --------------------- Receive Ports - RX Equalizer Ports -------------------
      gt0_rxdfelpmreset_in            =>      gt0_rxdfelpmreset_in,
      gt0_rxmonitorout_out            =>      gt0_rxmonitorout_out,
      gt0_rxmonitorsel_in             =>      gt0_rxmonitorsel_in,
      --------------- Receive Ports - RX Fabric Output Control Ports -------------
      gt0_rxoutclkfabric_out          =>      gt0_rxoutclkfabric_out,
      ------------- Receive Ports - RX Initialization and Reset Ports ------------
      gt0_gtrxreset_in                =>      gt0_gtrxreset_in,
      gt0_rxpmareset_in               =>      gt0_rxpmareset_in,
      ------------------- Receive Ports - RX8B/10B Decoder Ports -----------------
      gt0_rxcharisk_out               =>      gt0_rxcharisk_out,
      -------------- Receive Ports -RX Initialization and Reset Ports ------------
      gt0_rxresetdone_out             =>      gt0_rxresetdone_out,
      --------------------- TX Initialization and Reset Ports --------------------
      gt0_gttxreset_in                =>      gt0_gttxreset_in,
      gt0_txuserrdy_in                =>      gt0_txuserrdy_in,
      ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
      gt0_txusrclk_in                 =>      gt0_txusrclk_i,
      gt0_txusrclk2_in                =>      gt0_txusrclk2_i,
      ------------------ Transmit Ports - TX Data Path interface -----------------
      gt0_txdata_in                   =>      gt0_txdata_in,
      ---------------- Transmit Ports - TX Driver and OOB signaling --------------
      gt0_gtxtxn_out                  =>      gt0_gtxtxn_out,
      gt0_gtxtxp_out                  =>      gt0_gtxtxp_out,
      ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
      gt0_txoutclk_out                =>      gt0_txoutclk_i,
      gt0_txoutclkfabric_out          =>      gt0_txoutclkfabric_out,
      gt0_txoutclkpcs_out             =>      gt0_txoutclkpcs_out,
      --------------------- Transmit Ports - TX Gearbox Ports --------------------
      gt0_txcharisk_in                =>      gt0_txcharisk_in,
      ------------- Transmit Ports - TX Initialization and Reset Ports -----------
      gt0_txresetdone_out             =>      gt0_txresetdone_out,



      gt0_qplloutclk_in    =>GT0_QPLLOUTCLK_OUT,
      gt0_qplloutrefclk_in =>GT0_QPLLOUTREFCLK_OUT
      );



end RTL;


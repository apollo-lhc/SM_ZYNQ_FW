ibert_top.vhd
sdsdssd

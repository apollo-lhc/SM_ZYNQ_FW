../rev1_xc7z035/top.vhd
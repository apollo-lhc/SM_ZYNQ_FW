module gf_add_4(op1, op2, res);

// -------------------------------------------------------------------------- //
// ------------- Triple Modular Redundancy Generator Directives ------------- //
// -------------------------------------------------------------------------- //
// tmrg do_not_touch
// -------------------------------------------------------------------------- //

	input      [3:0] op1; 
	input      [3:0] op2; 
	output     [3:0] res;

	assign res = op1 ^ op2;

endmodule

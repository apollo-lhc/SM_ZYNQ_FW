../rev2_xc7z035/top.vhd